module
C_GEN (J,K,F5);
input J,K;
output F5;
xor G1(F5,J,K);
endmodule
